module crc_two
	(
		input i_rst_n,
		input i_clk,

		input i_data,
		output o_code
	);

	reg r_code;

	reg r_d0;
	reg r_d1;
	reg r_d2;
	reg r_d3;



endmodule
